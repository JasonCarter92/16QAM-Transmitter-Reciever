module SUT(	
				input sys_clk,
				input sym_clk_ena,
				input sam_clk_ena,
				input SW;
				input [1:0] mapperIn,
				output reg [17:0] decisionVariable);
				
				

			
endmodule	

				