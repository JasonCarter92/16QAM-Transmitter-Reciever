module ErrorGen ();

endmodule
